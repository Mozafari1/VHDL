----------------------------------------------------------------------------------
-- Company: 
-- Engineer: KIRISAN & RAHMAT
-- 
-- Create Date: 15.10.2019 22:38:16
-- Design Name: 
-- Module Name: top_tb - arch
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 -- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
ENTITY top_tb IS
END top_tb;
 
ARCHITECTURE behavior of top_tb is 
 
    -- Component Declarations for the Units Under Test (UUT)
    COMPONENT top
	port(
			clk, rst: in std_logic;
			ob: out std_logic_vector(7 downto 0)
		);
    END COMPONENT;

   --Inputs
   signal clk,rst : std_logic := '0';
   --Outputs
   signal ob : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	--Unit Under Test (UUT)
   uut: top PORT MAP (
          clk => clk,
          rst => rst, 
          ob => ob

        );

   -- Clock process 
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_pro: process
   begin		
        rst <= '1';
        wait for clk_period*2;
		rst <= '0';	
		wait for clk_period*2000000000;

   end process;

END;

